// megafunction wizard: %ALTUFM_SPI%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTUFM_SPI 

// ============================================================
// File Name: spi.v
// Megafunction Name(s):
// 			ALTUFM_SPI
//
// Simulation Library Files(s):
// 			maxii
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.1 Build 243 01/31/2013 SP 1 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module spi (
	ncs,
	sck,
	si,
	so)/* synthesis synthesis_clearbox = 1 */;

	input	  ncs;
	input	  sck;
	input	  si;
	output	  so;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX II"
// Retrieval info: PRIVATE: OSC_PORT STRING "OFF"
// Retrieval info: CONSTANT: ACCESS_MODE STRING "READ_ONLY"
// Retrieval info: CONSTANT: BYTE_OF_PAGE_WRITE NUMERIC "8"
// Retrieval info: CONSTANT: CONFIG_MODE STRING "EXTENDED"
// Retrieval info: CONSTANT: ERASE_TIME NUMERIC "500000000"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX II"
// Retrieval info: CONSTANT: LPM_FILE STRING "/home/jiakai/document/original/thu/2013-spring/assignment/digit-circuit/blxlrsmb/gen/mem.mif"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altufm_spi"
// Retrieval info: CONSTANT: OSC_FREQUENCY NUMERIC "180000"
// Retrieval info: CONSTANT: PROGRAM_TIME NUMERIC "1600000"
// Retrieval info: CONSTANT: WIDTH_UFM_ADDRESS NUMERIC "9"
// Retrieval info: USED_PORT: ncs 0 0 0 0 INPUT NODEFVAL "ncs"
// Retrieval info: CONNECT: @ncs 0 0 0 0 ncs 0 0 0 0
// Retrieval info: USED_PORT: sck 0 0 0 0 INPUT NODEFVAL "sck"
// Retrieval info: CONNECT: @sck 0 0 0 0 sck 0 0 0 0
// Retrieval info: USED_PORT: si 0 0 0 0 INPUT NODEFVAL "si"
// Retrieval info: CONNECT: @si 0 0 0 0 si 0 0 0 0
// Retrieval info: USED_PORT: so 0 0 0 0 OUTPUT NODEFVAL "so"
// Retrieval info: CONNECT: so 0 0 0 0 @so 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL spi.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL spi.cmp TRUE TRUE
// Retrieval info: LIB_FILE: maxii
